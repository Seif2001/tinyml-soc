module i2s(
    input clk,
    input rst_n,
    output WS,
    output BCLK,
    input DIN,
);





endmodule